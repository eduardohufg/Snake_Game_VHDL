LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY VGA_CONTROLLER IS
	PORT(CLK, RST, START: IN STD_LOGIC;
			ENAB: OUT STD_LOGIC;
			HSYNC, VSYNC: OUT STD_LOGIC;
			FIL, COL: OUT STD_LOGIC_VECTOR (9 DOWNTO 0));
			
	END VGA_CONTROLLER;
	
	
ARCHITECTURE RTL OF VGA_CONTROLLER IS

	
	COMPONENT DIVFREQ2 IS
	port(
		clk, reset: in std_logic;
		F: OUT STD_logic);
		END COMPONENT DIVFREQ2;
		
		
	COMPONENT CONT800 IS
	PORT(CLK, RST: IN STD_LOGIC; --Bits de control
			O: OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
			ov: out std_LOGIC); --Over Flow del contador
	END COMPONENT CONT800;
	
	
	COMPONENT CONTMOD525 IS
	PORT(CLK, RST: IN STD_LOGIC; --Bits de control
			O: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)); --Over Flow del contador
	END COMPONENT CONTMOD525;
	
	COMPONENT MESTADOSVSYNC IS
   --	entradas de control, tiempos y salidas
	PORT ( RST, CLK, START: IN std_logic;
			 CUENTA    :  IN std_logic_vector(9 DOWNTO 0);
			 VSYNC: OUT STD_logic;
			 VA: OUT STD_logic);
		END COMPONENT MESTADOSVSYNC; 
	
	
	COMPONENT MESTADOSHSYNC IS
   --	entradas de control, tiempos y salidas
	PORT ( RST, CLK, START: IN std_logic;
			 CUENTA    :  IN std_logic_vector(9 DOWNTO 0);
			 HSYNC: OUT STD_logic;
			 VA: IN STD_logic;
			 ENA: OUT STD_logic;
			 CUENTAV: IN STD_logic_vector(9 DOWNTO 0));
		end COMPONENT MESTADOSHSYNC;
	
		
	SIGNAL CLK25MHZ: STD_LOGIC;
	SIGNAL CONTA800: STD_LOGIC_VECTOR (9 DOWNTO 0);
	SIGNAL CONT525: STD_LOGIC_VECTOR (9 DOWNTO 0);
	SIGNAL OV800: STD_LOGIC;
	SIGNAL VAC: STD_LOGIC;
		
		
	
	BEGIN
	
		I0: DIVFREQ2 PORT MAP (CLK, RST, CLK25MHZ);
		I1: CONT800 PORT MAP(CLK25MHZ, RST, CONTA800, OV800);
		I2: CONTMOD525 PORT MAP(OV800, RST, CONT525);
		I3: MESTADOSVSYNC PORT MAP(RST, CLK25MHZ, START, CONT525, VSYNC, VAC);
		I4: MESTADOSHSYNC PORT MAP(RST,CLK25MHZ, START,CONTA800, HSYNC, VAC, ENAB, CONT525);
		
		
	
		FIL<= CONT525;
		COL<= CONTA800;
		
	END RTL;
	


	